library ieee;
use ieee.std_logic_1164.all;

package globals is
	constant NBIT : integer := 32;
end globals;
